module ID_EX_reg
(

);

endmodule